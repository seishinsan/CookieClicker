1.0
2.5599999999999996
21.679999999999996
60.0
100.0
150.0