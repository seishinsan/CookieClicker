7.46
30.714266438417116
331.46147926398856
179.15903999999998
180.0
525.0